`timescale 1ns/1ps

module buffer(
  input  wire gi,
  output wire g
);

assign g = gi;

endmodule
